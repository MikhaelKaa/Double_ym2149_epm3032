`timescale 1ns/1ps
module EPM3032_YM2149x2 (
input a0, a1, a2, a14, a15,
input cpu_clock, m1, iorq, wr, int, 
input reset,  
input d_0, d_3, d_4, d_5, d_6, d_7,  
//input d7_alt,
input dos,
output covox, 

output bc1, 
output bdir, 
output ym_clock, 
output ym_0, ym_1,
output beeper,
output tapeout,
output ioge_c,
output test
);

// Для тактирования звукового генератора 3.5.
//assign ym_clock = cpu_clock;


// Для тактирования звукового генератора при изменении частоты 7\3.5.
reg [14:0] clk_div_cnt = 0;
reg clk_div2 = 0; 
reg clk_detect_70m = 0;

always @(negedge cpu_clock) begin
	clk_div2 = ~clk_div2;
	if(int) begin 
		clk_div_cnt = clk_div_cnt + 1;
	end
	else begin 
		if(clk_div_cnt[14]) begin
			clk_div_cnt <= 0;
			clk_detect_70m = clk_div_cnt[14];
		end 
		else clk_div_cnt = 0;
	end
end	

/*always @(negedge int) begin
	clk_check7 = ~clk_check7;
	clk_detect_70m = clk_div_cnt[18];
end*/


assign ym_clock = (clk_detect_70m)?(clk_div2):(cpu_clock);


//assign test = clk_detect_70m;

// covox
assign covox = ~(a2 | iorq | wr | ~dos);

// Дешифрация звукового генератора.
wire   ssg 	= ~(a15 & (~(a1 | iorq)));
assign bc1  = ~(ssg | (~(a14 & m1)));
assign bdir = ~(ssg | wr);

// IORQGE
assign ioge_c = bc1 | bdir;

// Turbo Sound
reg  YM_select = 1'b0;
wire TS_bit_sel = ~(d_3 & d_4 & d_5 & d_6 & d_7 & bdir & bc1); 
//wire TS_bit_sel = ~(d_3 & d_4 & d_5 & d_6 & d7_alt & bdir & bc1); 
always @(negedge TS_bit_sel or negedge reset) begin
	if(~reset) 	YM_select = 1'b0;
	else 			YM_select = d_0;
end
assign ym_0 = ~YM_select;
assign ym_1 = ~ym_0;



// Дешифрация бипера и tapeout. Аналогично пентагоновской схеме.

// d7 on 26 pin
reg pre_beeper = 0;
reg pre_tapeout = 0;
always @(negedge wr) begin
	if( ~( iorq | a0) ) pre_beeper  = d_4;
	if( ~( iorq | a0) ) pre_tapeout = d_3;
end
assign beeper = pre_beeper;
assign tapeout = pre_tapeout;
//assign tapeout = dos;



/*
// d7 on 33 pin
reg pre_beeper;
reg pre_tapeout;
always @(negedge cpu_clock) begin
	if( ~(iorq | wr | a0) ) pre_beeper  = d[4];
	if( ~(iorq | wr | a0) ) pre_tapeout = d[3];
end

assign beeper = pre_beeper;
assign tapeout =  pre_tapeout;*/



//assign beeper = 1'bz;
//assign tapeout = 1'bz;

endmodule